module d_ff(D,clock,Q,Qbar)
input D,clock;
reg Q,Qbar;
assign ;
end module 