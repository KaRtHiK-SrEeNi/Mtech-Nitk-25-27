module and_stc(Y,A,B);
    input A,B;
    output Y;
    and gate( Y, A, B );
endmodule